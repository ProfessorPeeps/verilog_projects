/********************************************************************
 ***														   	  ***
 *** EE 526 L Experiment #10		   Juan Silva, Spring 2019    ***
 *** 														   	  ***
 *** Modeling a Sequencer Controller							  ***
 ********************************************************************
 *** Filename: phaser.sv		 	Created By Juan Silva 4/11/19 ***
 ***														   	  ***
 ********************************************************************
 ********************************************************************/
 `timescale 1 ns / 1 ns
 
 module RISCY(CLK, RST, IO);
 
output IO;
input CLK, RST;
 
//Instantiate necessary modules

	/*
	sequencer 		seq1(
	top_counter 	cnt1(
	scale_mux 		MUX1(
	alu				ALU1(
	AASD			aasd1(
	*/
	
	
endmodule