/********************************************************************
 ***														   	  ***
 *** EE 526 L Experiment #10		   Juan Silva, Spring 2019    ***
 *** 														   	  ***
 *** Modeling a Sequencer Controller							  ***
 ********************************************************************
 *** Filename: sequencer.sv		 	Created By Juan Silva 4/11/19 ***
 ***														   	  ***
 ********************************************************************
 *** 
 ********************************************************************/
 
`timescale 1 ns / 1 ns
 
module  RISCY(CLK, RST, IO);

input CLK, RST;
input [7:0] IO;

endmodule
	
